`ifndef _blob_vh_
`define _blob_vh_

`define BLOB_WIDTH   75

`define VALID        0:0
`define EQ_IND       9:1
`define COUNT        29:10
`define MIN_I        40:30
`define MAX_I        51:41
`define MIN_J        62:52
`define MAX_J        73:63
`define FIRST_CLEAR  74:74

`endif  //_blob_vh_

